// FILE NAME: SRAM_TB.v
// TYPE: module_TB
// AUTHOR: Ahmed Gomaa
// AUTHOR’S EMAIL:ahmed.gomaa.work150@gmail.com
//---------------------------------------------------------------------
// PURPOSE: Digital Design Test Bench Project
//---------------------------------------------------------------------
// KEYWORDS: SRAM Test Bench
//---------------------------------------------------------------------
// Copyright 2024, Ahmed Gomaa, All rights reserved.
//---------------------------------------------------------------------

////////////////////////////////////////////////////////
//////////////// Module Difinition ///////////////////// 
////////////////////////////////////////////////////////

module SRAM_TB ();


////////////////////////////////////////////////////////
/////////////////// DUT Signals //////////////////////// 
////////////////////////////////////////////////////////

reg                               CLK   ;     // clock domain
reg          [ 3 : 0  ]           ADDR  ;     // address
reg          [ 7  : 0 ]           WDATA ;     // write data
reg                               WREN  ;     // write enable
wire         [ 7  : 0 ]           RDATA ;      // read data


////////////////////////////////////////////////////////
////////////////// initial block /////////////////////// 
////////////////////////////////////////////////////////

initial 
begin
    $dumpfile("SRAM.vcd") ;       // Save Waveform
    $dumpvars;
    CLK  = 0  ;
    WREN = 0 ;   ADDR = 4'b 0000 ;   WDATA = 8'b 0000_0000 ;  #10
    WREN = 1 ;   ADDR = 4'b 0001 ;   WDATA = 8'b 1010_1010 ;  #10
    WREN = 0 ;   ADDR = 4'b 0001 ;   WDATA = 8'b 0000_0000 ;  #10 $finish ;
end


////////////////////////////////////////////////////////
////////////////// Clock Generator  ////////////////////
////////////////////////////////////////////////////////

always    #5       CLK = ~ CLK  ;

////////////////////////////////////////////////////////
/////////////////// DUT Instantation ///////////////////
////////////////////////////////////////////////////////

SRAM DUT (    CLK  ,    ADDR  ,    WDATA  ,    WREN  ,    RDATA ) ;

endmodule



